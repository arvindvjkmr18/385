module position_subsystem(

	// Input timing:
	input logic				CLOCK_50,		// Master data clock
	input logic				PS2_CLK,			// PS2 Protocol clock
	
	// Input control:
	input logic				RESET_H,			// Reset command (active high)
	input logic				RUN_POS_UPDATE,// Control signal from system core FSM
	
	// Input data:
	input logic 			PS2_DAT,
	input logic	[1:0] 	SPRITE_ID,		// from Entity File
	input logic [8:0]		TARGET_X,		// entity's stored x,y coords
	input logic [8:0]		TARGET_Y,
	input logic [2:0]		STOP_ADDRESS,	
	
	// Output control:
	output logic			POS_UPDATE_DONE,// Communication back to system core FSM
	output logic			GAME_OVER,		// Indication of game over event
	output logic			YOU_WIN,
	output logic			WE_reg,
	
	// Output data:
	output logic [1:0]	ADDRESS,			// Entity file address
	output logic [1:0]	SPRITE_ID_reg,	// Sprite ID Code to assign for entity at address
	output logic [8:0]	TARGET_X_reg,	// Updated x,y coords...
	output logic [8:0]	TARGET_Y_reg,
	
	output logic [6:0]	HEX0, HEX1
	
	//output logic COLLISION, POS_CTRL_DEBUG

);

	// Internal wires:
	logic collision_done, get_input, trigger_ai, buffer_load, run_collision, game_over_flag, you_win_flag;
	logic [1:0] addr_mux_sel;
   logic	buf_mux_sel;
	logic [1:0] fsm_addr, collision_addr, collision_mux_addr, buf_mux_addr, buf_addr;
	logic [1:0] buf_mux_code, buf_code, collision_code, collision_mux_code;
	logic [8:0] buf_mux_x, buf_mux_y, buf_x, buf_y, hero_x, hero_y, enemy_x, enemy_y, collision_x, collision_y, collision_mux_x, collision_mux_y;
	
	// Other assignments:
	assign SPRITE_ID_reg = buf_code;
	assign TARGET_X_reg = buf_x;
	assign TARGET_Y_reg = buf_y;
	
	
	// Controller for position subsystem
	positionController FSM(
	
		.CLOCK_50,
		.RESET_H,
		.RUN_POS_UPDATE,
		.COLLISION_DONE(collision_done),
		.GAME_OVER_FLAG(game_over_flag),
		.YOU_WIN_FLAG(you_win_flag),
		.STOP_ADDRESS,
		.ID_CODE(SPRITE_ID),
		.POS_UPDATE_DONE,
		.GAME_OVER,
		.YOU_WIN,
		.GET_INPUT(get_input),
		.TRIGGER_AI(trigger_ai),
		.BUFFER_LOAD(buffer_load),
		.RUN_COLLISION(run_collision),
		.ADDR_MUX_SEL(addr_mux_sel),
		.BUF_MUX_SEL(buf_mux_sel),
		.WE_reg,
		.ADDRESS(fsm_addr)
	
	);
	
	// Controls access to the ADDRESS port (to the Entity File)
	addr_MUX addr_out_control(
	
		.SEL(addr_mux_sel),			// Select signal from FSM
		.ADDR_A(fsm_addr),	// Addr from Detect Collision module
		.ADDR_B(buf_addr),			// Addr from position buffer
		.ADDR_C(collision_addr),
		.ADDR_OUT(ADDRESS)			// Output to ADDRESS output port
	
	);

	// Controls access to the local entity buffer
	opcode_MUX pos_buf_mux(
	
		.SEL(buf_mux_sel),
		// Entity File input
		.ADDR_A(fsm_addr),		// Address generated by FSM
		.ID_CODE_A(SPRITE_ID),
		.X_A(TARGET_X),
		.Y_A(TARGET_Y),
		// Collision detection input
		.ADDR_B(collision_mux_addr),
		.ID_CODE_B(collision_code),
		.X_B(collision_x),
		.Y_B(collision_y),
		// Output
		.ADDR_OUT(buf_mux_addr),
		.ID_CODE_OUT(buf_mux_code),
		.X_OUT(buf_mux_x),
		.Y_OUT(buf_mux_y)
	
	);
	
	// Stores local copy of sprite opcode data for updating
	position_buffer entity_buffer(
	
		.CLOCK_50,
	
		.BUFFER_LOAD(buffer_load),

		.ADDR_IN(buf_mux_addr),
		.ID_CODE_IN(buf_mux_code),
		.X_IN(buf_mux_x),
		.Y_IN(buf_mux_y),
	
		.ADDR_OUT(buf_addr),
		.ID_CODE_OUT(buf_code),
		.X_OUT(buf_x),
		.Y_OUT(buf_y)
	
	);

	// Captures user input from PS/2 KB and applies it to new position (i.e. player motion)
	user_control_system player(
		
		// Input timing signals:
		.CLOCK_50,
		.PS2_CLK,
		.RESET_H,
	
		// Input control signals:
		.GET_INPUT(get_input),	// From module's FSM
	
		// Input data
		.PS2_DAT,					// From PS2 keyboard
		.CURR_POS_X(buf_x),		// Hero x,y from entity file
		.CURR_POS_Y(buf_y),
	
		// Output data
		.HERO_NEW_X(hero_x),		// New x,y position to entity file
		.HERO_NEW_Y(hero_y),

		// For visual keyboard input verification
		.HEX0, 
		.HEX1
	
	);
	
	// References last player position and derives new AI postion (i.e. AI motion)
	ai_control_system enemy(
	
		.CLOCK_50,
		.RESET_H,
		
		.RUN_AI(trigger_ai),
		.GET_PLAYER_POS(get_input),
		.PLAYER_X(TARGET_X),
		.PLAYER_Y(TARGET_Y),
		
		.TARGET_X(buf_x),
		.TARGET_Y(buf_y),
		
		.NEW_ENEMY_X(enemy_x),
		.NEW_ENEMY_Y(enemy_y)
	
	);
	
	// Controls access to the collision detection routine circuits
	opcode_MUX collision_mux(
	
		.SEL(buf_code[0]),		// This will need to be changed as more sprite IDs are added...
		// Entity File input
		.ADDR_A(buf_addr),		// Address generated by FSM
		.ID_CODE_A(buf_code),
		.X_A(hero_x),
		.Y_A(hero_y),
		// Collision detection input
		.ADDR_B(buf_addr),
		.ID_CODE_B(buf_code),
		.X_B(enemy_x),
		.Y_B(enemy_y),
		// Output
		.ADDR_OUT(collision_mux_addr),
		.ID_CODE_OUT(collision_mux_code),
		.X_OUT(collision_mux_x),
		.Y_OUT(collision_mux_y)
	
	);
	
	// Collision detection routine circuits; confirms new position is valid
	detect_collision dc_comp(
	
		// Input timing
		.CLOCK_50,
	
	// Input control
		.RUN_COLLISION(run_collision),
		//.PLAYER_MOTION,						// Flag for whether player or monster is being checked.
		.STOP_ADDRESS,
	
	// Input data
		.MOVER_ID(collision_mux_code),
		.OLD_X(buf_x),							// Moving entity old x,y coord
		.OLD_Y(buf_y),
		.NEW_X(collision_mux_x),			// Moving entity new x,y coord
		.NEW_Y(collision_mux_y),
	
		.OBJ_ID(SPRITE_ID),					// Obstacle ID code
		.OBJ_X(TARGET_X),						// Obstacle obj x,y coord
		.OBJ_Y(TARGET_Y),
	
	// Output control
		.COLLISION_DONE(collision_done),// Command to position subsys FSM
		.GAME_OVER_FLAG(game_over_flag),// Game over condition flag
		.YOU_WIN_FLAG(you_win_flag),	  // i win
		
	// Output data
		.ADDRESS(collision_addr),			// Address for reading from entity file
		.ID_CODE(collision_code),			// Sprite ID code of collision-checked entity
		.FINAL_X(collision_x),				// Collision-checked x,y coord for moving entity
		.FINAL_Y(collision_y)
		
	);	

endmodule